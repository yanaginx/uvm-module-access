// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: arith_monitor.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Thu Nov 10 00:04:59 2022
//=============================================================================
// Description: Monitor for arith
//=============================================================================

`ifndef ARITH_MONITOR_SV
`define ARITH_MONITOR_SV

// You can insert code here by setting monitor_inc_before_class in file arith.tpl

class arith_monitor extends uvm_monitor;

  `uvm_component_utils(arith_monitor)

  virtual arith_if vif;

  arith_config     m_config;

  uvm_analysis_port #(trans) analysis_port;

  trans m_trans;

  extern function new(string name, uvm_component parent);

  // Methods run_phase, and do_mon generated by setting monitor_inc in file arith.tpl
  extern task run_phase(uvm_phase phase);
  extern task do_mon();

  // You can insert code here by setting monitor_inc_inside_class in file arith.tpl

endclass : arith_monitor 


function arith_monitor::new(string name, uvm_component parent);
  super.new(name, parent);
  analysis_port = new("analysis_port", this);
endfunction : new


task arith_monitor::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  m_trans = trans::type_id::create("m_trans");
  do_mon();
endtask : run_phase


// Start of inlined include file generated_tb/tb/include/arith_monitor_inc.sv
task arith_monitor::do_mon;
  forever @(vif.F)
  begin
    m_trans.input1 = vif.A;
    m_trans.input2 = vif.B;
    m_trans.sum    = vif.F;
    analysis_port.write(m_trans);
    `uvm_info(get_type_name(), 
                $sformatf("%0d + %0d = %0d", 
                            vif.A,
                            vif.B,
                            vif.F),
                UVM_MEDIUM) 
  end
endtask
// End of inlined include file

// You can insert code here by setting monitor_inc_after_class in file arith.tpl

`endif // ARITH_MONITOR_SV

